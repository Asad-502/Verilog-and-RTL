
module statemachine1(x,y,clock,reset);
input x,clock,reset;
output y;
reg y;
reg [1:0]prstate,nxtstate;
parameter s0=2'b00 , s1=2'


endmodule
